-- Code your testbench here
library IEEE;
use IEEE.std_logic_1164.all;

entity Testbench is  
end Testbench; 